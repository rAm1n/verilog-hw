module bcd_greey(a,b,c,d,in);
    input [3:0] in ;
    output a,b,c,d ;
    assign {a,b,c,d} = (in == 4'b 0000) ? 4'b 0000 :
			 (in == 4'b 0001) ? 4'b 0001 :
			 (in == 4'b 0010) ? 4'b 0011 :
			 (in == 4'b 0011) ? 4'b 0010 :
			 (in == 4'b 0100) ? 4'b 0110 :
			 (in == 4'b 0101) ? 4'b 0111 :
			 (in == 4'b 0110) ? 4'b 0101 :
			 (in == 4'b 0111) ? 4'b 0100 :
			 (in == 4'b 1000) ? 4'b 1100 :
			 (in == 4'b 1001) ? 4'b 1101 :
			 (in == 4'b 1010) ? 4'b 1111 :
			 (in == 4'b 1011) ? 4'b 1110 :
			 (in == 4'b 1100) ? 4'b 1010 :
			 (in == 4'b 1101) ? 4'b 1011 :
			 (in == 4'b 1110) ? 4'b 1001 :
			 (in == 4'b 1111) ? 4'b 1000 : 4'b0000 ;
endmodule
